* C:\LTspice\examples\Educational\waveout.cir
.end
