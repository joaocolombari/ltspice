* U:\LTspice\examples\jigs\1009.asc
V1 N001 0 0
R1 N001 OUT 3.6K
XU1 OUT 0 N002 LT1009
R2 OUT N002 {10K*(1-x)}
R3 N002 0 {10K*x}
.dc TEMP -55 125 .1
.step param x .4 .6 .1
.lib LTC3.lib
.backanno
.end
